module moore (
input clk, reset, x,        
output reg z              
);
parameter S0 = 3'b000,  
          S1 = 3'b001,  
          S2 = 3'b010,  
          S3 = 3'b011,  
          S4 = 3'b100;  
reg [2:0] state, next_state;
always @(posedge clk or posedge reset) 
begin
if (reset)
state <= S0;
else
state <= next_state;
end
always @(*) begin
case (state)
 S0: next_state = (x) ? S1 : S0;
 S1: next_state = (x) ? S1 : S2;
 S2: next_state = (x) ? S3 : S0;
 S3: next_state = (x) ? S4 : S2;
 S4: next_state = (x) ? S1 : S2;
 default: next_state = S0;
endcase
end
always @(*) 
begin
case (state)
 S4: z = 1'b1;
default: z = 1'b0;
endcase
end

endmodule

